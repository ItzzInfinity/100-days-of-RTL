`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Anjan Prasad
// Create Date: 11/24/2024 05:19:14 AM
// Module Name: half_adder
//////////////////////////////////////////////////////////////////////////////////

module half_adder(
	input a,b,
	output sum,carry
	);
    assign sum=a^b;
    assign carry=a&b;
endmodule