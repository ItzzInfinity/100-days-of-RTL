
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Anjan Prasad
// Create Date: 10/23/2024 06:11:25 AM
// Module Name: mux_4_to_1
//////////////////////////////////////////////////////////////////////////////////


module mux_4_to_1(
    input [3:0]a,
    input [1:0] sel,
    output y);
    
        assign y = a[sel];

endmodule
