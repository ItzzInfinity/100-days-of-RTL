
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Anjan Prasad
// Create Date: 10/22/2024 06:16:32 AM
// Module Name: demux_1_to_2
//////////////////////////////////////////////////////////////////////////////////

module demux_1_to_2(
    input sel,
    input i,
    output y0, y1
    );    
    assign {y0,y1} = sel?{1'b0,i}: {i,1'b0};
endmodule